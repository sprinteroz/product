.TITLE Full Wave Rectifier
V1 3 2 SIN(0.0 208.0 159.15)
RL 1 GND 1k
//Diode D1
D1 GND 3 dmod_d1 area=1 ic=0.0
.MODEL dmod_d1 D (level=1)
//Diode D3
D3 2 1 dmod_d3 area=1 ic=0.0
.MODEL dmod_d3 D (level=1)
//Diode D4
D4 3 1 dmod_d4 area=1 ic=0.0
.MODEL dmod_d4 D (level=1)
//Diode D2
D2 GND 2 dmod_d2 area=1 ic=0.0
.MODEL dmod_d2 D (level=1)
.TRAN 50µ 25m
.PRINT TRAN v(1) @Rl[i]
.END