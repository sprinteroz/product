.TITLE Bipolar Amplifier
Vin in GND SIN(0.0 1m 500.0)
Vcc cc GND 5.0
R1 cc intb 68k
R3 cc intc 10k
Cin in intb 10µ
Cout intc out 10µ
RLoad out GND 100k
R2 intb GND 10k
Q1 intc intb GND qmod_q1
.MODEL qmod_q1 NPN level=1 vaf=73.4 is=7.590f vjc=650m rb=100.0
+ vje=650m rc=250m re=500m rbm=10.0 bf=480.0 br=5.0 irb=100µ
+ mje=550m vtf=3.0 tf=426p isc=200f ise=3.278f tr=150n ikf=96.200m
+ ikr=30m itf=600m nc=1.2 ne=1.2665 cjc=6.330p cje=12.500p xtf=20.0
.TRAN 10µ 10m
.PRINT TRAN v(out) v(in)
.END