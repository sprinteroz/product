.TITLE RC AC
R1 GND 1 5k
C1 1 GND 20n IC=5.0
.TRAN 5µ 1m UIC
.PRINT TRAN v(1)
.END